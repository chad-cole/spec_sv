package database_pkg; 

`include "macros.svh"
`include "factory.sv"
`include "file_string_tasks.sv"
`include "database.sv"

endpackage : database_pkg
